// instruction memory
module scinstmem (pc, inst);


endmodule
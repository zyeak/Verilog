// data memory
module scdatamem (clk, mem_out, data, alu_out, wmen);


endmodule